test AMP_IDC_CurrentBias

.LIB '../models/sky130.lib.spice'tt
.INCLUDE AMP_CurrentBias.cir
.INCLUDE CurrentBias.cir


V1 VSS 0 dc=0V
V0 VDD_SOURCE 0 dc=1.8V
VMEAS VDD_SOURCE VDD 0

VIN Vinn 0 dc=0.9V
VIP Vinp 0 dc=0.9V

XI1 Vinp Vinn VDD VSS Vout AMP_CurrentBias
C1 VOUT 0 2E-12

.CONTROL
set units=degrees
run
op
print i(vmeas) >Idc.txt


.ENDC
.END
