test AMP_PSRR

.LIB '/mnt/c/llm/package/models/sky130.lib.spice'tt
.INCLUDE /mnt/c/llm/LLM4AMP/agent/sim_src/AMP.cir
.TEMP 25.0

V1 VSS 0 dc=0V
V0 VDD 0 dc=1.8V ac=1
VIP Vinp 0 dc=0.9V

XI1 Vinp Vout VDD VSS Vout AMP
C1 VOUT 0 2E-12

.control
set units = degrees
run

compose ac_pts start=1 stop=1e6 dec=10
let freq_pts = ac_pts

ac dec 10 1 1Meg
meas ac vdd_gain find vdb(VOUT) at=1e3Hz
let vdd_gain1 = -vdd_gain
echo "$&vdd_gain1" > /mnt/c/llm/LLM4AMP/agent/sim_result/ttPSRR_results.txt
plot vdb(VOUT)

quit
.ENDC
.END
