test AMP_IDC_CurrentBias

.LIB '/root/submission/final_netlist2/models/sky130.lib.spice'ss
.INCLUDE /root/submission/final_netlist2/AMP.cir
.INCLUDE /root/submission/final_netlist2/CurrentBias.cir


V1 VSS 0 dc=0V
V0 VDD_SOURCE 0 dc=1.8V
VMEAS VDD_SOURCE VDD 0

VIN Vinn 0 dc=0.9V
VIP Vinp 0 dc=0.9V

XI1 Vinp Vinn VDD VSS Vout AMP
C1 VOUT 0 2E-12

.CONTROL
set units=degrees
run
op
print i(vmeas) >SS_Idc.txt


.ENDC
.END
