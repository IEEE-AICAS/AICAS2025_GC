.subckt CurrentBias Ibias VDD VDD2 VSS

.param W12 = 8      	    mult_12 = 1  		    L12 = 1.0
.param W34 = 8    	    mult_34 = 1   			L34 = 1.0
.param W5_6_7 = 2.5         L5_6_7 = 1


XM1 net1 net2 net0 VSS sky130_fd_pr__nfet_01v8 L=L12 W=W12 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=40 m=40

XM2 net2 net2 VSS VSS sky130_fd_pr__nfet_01v8 L=L12 W=W12 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=mult_12 m=mult_12 

XM3 net3 net4 net1 VSS sky130_fd_pr__nfet_01v8 L=L34 W=W34 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=mult_34 m=mult_34 

XM4 net4 net4 net2 VSS sky130_fd_pr__nfet_01v8 L=L34 W=W34 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=mult_34 m=mult_34

XM5 net3 net3 VDD VDD sky130_fd_pr__pfet_01v8 L=L5_6_7 W=W5_6_7 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1

XM6 net4 net3 VDD VDD sky130_fd_pr__pfet_01v8 L=L5_6_7 W=W5_6_7 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1 

XM7 net5 net3 VDD2 VDD2 sky130_fd_pr__pfet_01v8 L=L5_6_7 W=W5_6_7 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1

XM8 net5 net5 Ibias VSS sky130_fd_pr__nfet_01v8 L=L34 W=W34 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=mult_34 m=mult_34


R0 net0 VSS 10K
C1 net0 VSS 0.01p m=1
C2 net2 VSS 0.15p m=1
.ends CurrentBias