test AMP_IDC

.LIB '/mnt/c/llm/package/models/sky130.lib.spice'tt
.INCLUDE /mnt/c/llm/LLM4AMP/agent/sim_src/AMP.cir


V1 VSS 0 dc=0V
V0 VDD_SOURCE 0 dc=1.8V
VMEAS VDD_SOURCE VDD 0

VIN Vinn 0 dc=0.9V
VIP Vinp 0 dc=0.9V

XI1 Vinp Vinn VDD VSS Vout AMP
C1 VOUT 0 2E-12

.CONTROL
set units=degrees
run
op


print @m.xi1.xm8.msky130_fd_pr__nfet_01v8[id]
print i(vmeas)

let result = @r.xi1.r2[i]
echo "$&result" > /mnt/c/llm/LLM4AMP/agent/sim_result/tt_I0_results.txt


quit
.ENDC
.END
