test AMP_AC_CurrentBias

.LIB '/root/submission/final_netlist2/models/sky130.lib.spice'sf
.INCLUDE /root/submission/final_netlist2/AMP.cir
.INCLUDE /root/submission/final_netlist2/CurrentBias.cir
.TEMP 25.0


V1 VSS 0 dc=0V
V0 VDD 0 dc=1.8V
VIN Vinn 0 dc=0.9V ac=-0.5V
VIP Vinp 0 dc=0.9V ac=0.5V

XI1 Vinp Vinn VDD VSS Vout AMP
C1 Vout 0 2E-12

.ac dec 100 1Hz 1000MegHz
.print ac vdb(Vout)
.print ac vp(Vout)

.CONTROL
set units = degrees
run

compose ac_pts start=1 stop=1e9 dec=100
let freq_pts = ac_pts


meas ac gain_max find vdb(Vout) at=1Hz
meas ac gbw when vdb(Vout)=0
meas ac phase_val find vp(Vout) when vdb(Vout)=0
let phase_margin = 180 + phase_val


echo "Gain: $&gain_max" > SF_AC_results.txt
echo "GBW: $&gbw" >> SF_AC_results.txt
echo "PM: $&phase_margin" >> SF_AC_results.txt

.ENDC
.END
